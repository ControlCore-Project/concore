`timescale 1ns/100ps

module funcRom(romout,zH);
	output [11:0] romout;
	input [7:0] zH;
	reg [11:0] romout;
	always @(zH)
		begin
			case(zH)
1 :romout = 2;
2 :romout = 2;
3 :romout = 2;
4 :romout = 2;
5 :romout = 2;
6 :romout = 2;
7 :romout = 2;
8 :romout = 2;
9 :romout = 2;
10 :romout = 2;
11 :romout = 2;
12 :romout = 2;
13 :romout = 2;
14 :romout = 2;
15 :romout = 2;
16 :romout = 2;
17 :romout = 2;
18 :romout = 2;
19 :romout = 2;
20 :romout = 2;
21 :romout = 2;
22 :romout = 2;
23 :romout = 2;
24 :romout = 2;
25 :romout = 2;
26 :romout = 2;
27 :romout = 2;
28 :romout = 2;
29 :romout = 2;
30 :romout = 2;
31 :romout = 2;
32 :romout = 2;
33 :romout = 2;
34 :romout = 2;
35 :romout = 2;
36 :romout = 2;
37 :romout = 2;
38 :romout = 2;
39 :romout = 2;
40 :romout = 2;
41 :romout = 2;
42 :romout = 2;
43 :romout = 2;
44 :romout = 2;
45 :romout = 2;
46 :romout = 2;
47 :romout = 2;
48 :romout = 2;
49 :romout = 2;
50 :romout = 2;
51 :romout = 2;
52 :romout = 2;
53 :romout = 2;
54 :romout = 2;
55 :romout = 2;
56 :romout = 2;
57 :romout = 2;
58 :romout = 2;
59 :romout = 2;
60 :romout = 2;
61 :romout = 2;
62 :romout = 2;
63 :romout = 2;
64 :romout = 2;
65 :romout = 2;
66 :romout = 2;
67 :romout = 2;
68 :romout = 2;
69 :romout = 2;
70 :romout = 2;
71 :romout = 2;
72 :romout = 2;
73 :romout = 2;
74 :romout = 2;
75 :romout = 2;
76 :romout = 2;
77 :romout = 2;
78 :romout = 2;
79 :romout = 2;
80 :romout = 2;
81 :romout = 2;
82 :romout = 2;
83 :romout = 2;
84 :romout = 2;
85 :romout = 2;
86 :romout = 2;
87 :romout = 2;
88 :romout = 2;
89 :romout = 2;
90 :romout = 2;
91 :romout = 2;
92 :romout = 2;
93 :romout = 2;
94 :romout = 2;
95 :romout = 2;
96 :romout = 2;
97 :romout = 2;
98 :romout = 2;
99 :romout = 2;
100 :romout = 2;
101 :romout = 2;
102 :romout = 2;
103 :romout = 2;
104 :romout = 2;
105 :romout = 2;
106 :romout = 2;
107 :romout = 2;
108 :romout = 2;
109 :romout = 2;
110 :romout = 2;
111 :romout = 2;
112 :romout = 2;
113 :romout = 2;
114 :romout = 2;
115 :romout = 2;
116 :romout = 2;
117 :romout = 2;
118 :romout = 2;
119 :romout = 2;
120 :romout = 2;
121 :romout = 2;
122 :romout = 2;
123 :romout = 2;
124 :romout = 2;
125 :romout = 2;
126 :romout = 2;
127 :romout = 2;
128 :romout = 2;
129 :romout = 2;
130 :romout = 2;
131 :romout = 2;
132 :romout = 2;
133 :romout = 2;
134 :romout = 2;
135 :romout = 2;
136 :romout = 2;
137 :romout = 2;
138 :romout = 2;
139 :romout = 2;
140 :romout = 2;
141 :romout = 2;
142 :romout = 2;
143 :romout = 2;
144 :romout = 2;
145 :romout = 2;
146 :romout = 2;
147 :romout = 2;
148 :romout = 2;
149 :romout = 2;
150 :romout = 2;
151 :romout = 2;
152 :romout = 2;
153 :romout = 2;
154 :romout = 2;
155 :romout = 2;
156 :romout = 2;
157 :romout = 2;
158 :romout = 2;
159 :romout = 2;
160 :romout = 2;
161 :romout = 2;
162 :romout = 2;
163 :romout = 2;
164 :romout = 3;
165 :romout = 3;
166 :romout = 3;
167 :romout = 3;
168 :romout = 3;
169 :romout = 3;
170 :romout = 3;
171 :romout = 3;
172 :romout = 4;
173 :romout = 4;
174 :romout = 4;
175 :romout = 4;
176 :romout = 4;
177 :romout = 5;
178 :romout = 5;
179 :romout = 5;
180 :romout = 6;
181 :romout = 6;
182 :romout = 6;
183 :romout = 7;
184 :romout = 7;
185 :romout = 8;
186 :romout = 8;
187 :romout = 9;
188 :romout = 10;
189 :romout = 10;
190 :romout = 11;
191 :romout = 12;
192 :romout = 13;
193 :romout = 14;
194 :romout = 15;
195 :romout = 16;
196 :romout = 18;
197 :romout = 19;
198 :romout = 21;
199 :romout = 23;
200 :romout = 24;
201 :romout = 27;
202 :romout = 29;
203 :romout = 31;
204 :romout = 34;
205 :romout = 37;
206 :romout = 40;
207 :romout = 44;
208 :romout = 47;
209 :romout = 51;
210 :romout = 56;
211 :romout = 61;
212 :romout = 66;
213 :romout = 72;
214 :romout = 78;
215 :romout = 85;
216 :romout = 92;
217 :romout = 101;
218 :romout = 109;
219 :romout = 119;
220 :romout = 129;
221 :romout = 141;
222 :romout = 153;
223 :romout = 166;
224 :romout = 181;
225 :romout = 196;
226 :romout = 213;
227 :romout = 232;
228 :romout = 252;
229 :romout = 273;
230 :romout = 297;
231 :romout = 322;
232 :romout = 350;
233 :romout = 379;
234 :romout = 411;
235 :romout = 445;
236 :romout = 482;
237 :romout = 522;
238 :romout = 565;
239 :romout = 611;
240 :romout = 661;
241 :romout = 714;
242 :romout = 771;
243 :romout = 831;
244 :romout = 896;
245 :romout = 965;
246 :romout = 1038;
247 :romout = 1117;
248 :romout = 1200;
249 :romout = 1287;
250 :romout = 1380;
251 :romout = 1478;
252 :romout = 1582;
253 :romout = 1690;
254 :romout = 1805;
255 :romout = 1924;
0 : romout =2;
//0 :romout = 2050;
endcase
end
endmodule
module slopeRom(romout,zH);
	output [6:0] romout;
	input [7:0] zH;
	reg [6:0] romout;
	always @(zH)
		begin
			case(zH)
0 : romout=0;
255 : romout=119;
254 : romout=114;
253 : romout=108;
252 : romout=103;
251 : romout=98;
250 : romout=92;
249 : romout=87;
248 : romout=82;
247 : romout=78;
246 : romout=73;
245 : romout=69;
244 : romout=64;
243 : romout=60;
242 : romout=56;
241 : romout=53;
240 : romout=49;
239 : romout=46;
238 : romout=42;
237 : romout=39;
236 : romout=37;
235 : romout=34;
234 : romout=31;
233 : romout=29;
232 : romout=27;
231 : romout=25;
230 : romout=23;
229 : romout=21;
228 : romout=19;
227 : romout=18;
226 : romout=17;
225 : romout=15;
224 : romout=14;
223 : romout=13;
222 : romout=12;
221 : romout=11;
220 : romout=10;
219 : romout=9;
218 : romout=8;
217 : romout=8;
216 : romout=7;
215 : romout=6;
214 : romout=6;
213 : romout=5;
212 : romout=5;
211 : romout=4;
210 : romout=4;
209 : romout=4;
208 : romout=3;
207 : romout=3;
206 : romout=3;
205 : romout=2;
204 : romout=2;
203 : romout=2;
202 : romout=2;
201 : romout=2;
200 : romout=1;
199 : romout=1;
198 : romout=1;
197 : romout=1;
196 : romout=1;
195 : romout=1;
194 : romout=1;
193 : romout=1;
192 : romout=0;
191 : romout=0;
190 : romout=0;
189 : romout=0;
188 : romout=0;
187 : romout=0;
186 : romout=0;
185 : romout=0;
184 : romout=0;
183 : romout=0;
182 : romout=0;
181 : romout=0;
180 : romout=0;
179 : romout=0;
178 : romout=0;
177 : romout=0;
176 : romout=0;
175 : romout=0;
174 : romout=0;
173 : romout=0;
172 : romout=0;
171 : romout=0;
170 : romout=0;
169 : romout=0;
168 : romout=0;
167 : romout=0;
166 : romout=0;
165 : romout=0;
164 : romout=0;
163 : romout=0;
162 : romout=0;
161 : romout=0;
160 : romout=0;
159 : romout=0;
158 : romout=0;
157 : romout=0;
156 : romout=0;
155 : romout=0;
154 : romout=0;
153 : romout=0;
152 : romout=0;
151 : romout=0;
150 : romout=0;
149 : romout=0;
148 : romout=0;
147 : romout=0;
146 : romout=0;
145 : romout=0;
144 : romout=0;
143 : romout=0;
142 : romout=0;
141 : romout=0;
140 : romout=0;
139 : romout=0;
138 : romout=0;
137 : romout=0;
136 : romout=0;
135 : romout=0;
134 : romout=0;
133 : romout=0;
132 : romout=0;
131 : romout=0;
130 : romout=0;
129 : romout=0;
128 : romout=0;
127 : romout=0;
126 : romout=0;
125 : romout=0;
124 : romout=0;
123 : romout=0;
122 : romout=0;
121 : romout=0;
120 : romout=0;
119 : romout=0;
118 : romout=0;
117 : romout=0;
116 : romout=0;
115 : romout=0;
114 : romout=0;
113 : romout=0;
112 : romout=0;
111 : romout=0;
110 : romout=0;
109 : romout=0;
108 : romout=0;
107 : romout=0;
106 : romout=0;
105 : romout=0;
104 : romout=0;
103 : romout=0;
102 : romout=0;
101 : romout=0;
100 : romout=0;
99 : romout=0;
98 : romout=0;
97 : romout=0;
96 : romout=0;
95 : romout=0;
94 : romout=0;
93 : romout=0;
92 : romout=0;
91 : romout=0;
90 : romout=0;
89 : romout=0;
88 : romout=0;
87 : romout=0;
86 : romout=0;
85 : romout=0;
84 : romout=0;
83 : romout=0;
82 : romout=0;
81 : romout=0;
80 : romout=0;
79 : romout=0;
78 : romout=0;
77 : romout=0;
76 : romout=0;
75 : romout=0;
74 : romout=0;
73 : romout=0;
72 : romout=0;
71 : romout=0;
70 : romout=0;
69 : romout=0;
68 : romout=0;
67 : romout=0;
66 : romout=0;
65 : romout=0;
64 : romout=0;
63 : romout=0;
62 : romout=0;
61 : romout=0;
60 : romout=0;
59 : romout=0;
58 : romout=0;
57 : romout=0;
56 : romout=0;
55 : romout=0;
54 : romout=0;
53 : romout=0;
52 : romout=0;
51 : romout=0;
50 : romout=0;
49 : romout=0;
48 : romout=0;
47 : romout=0;
46 : romout=0;
45 : romout=0;
44 : romout=0;
43 : romout=0;
42 : romout=0;
41 : romout=0;
40 : romout=0;
39 : romout=0;
38 : romout=0;
37 : romout=0;
36 : romout=0;
35 : romout=0;
34 : romout=0;
33 : romout=0;
32 : romout=0;
31 : romout=0;
30 : romout=0;
29 : romout=0;
28 : romout=0;
27 : romout=0;
26 : romout=0;
25 : romout=0;
24 : romout=0;
23 : romout=0;
22 : romout=0;
21 : romout=0;
20 : romout=0;
19 : romout=0;
18 : romout=0;
17 : romout=0;
16 : romout=0;
15 : romout=0;
14 : romout=0;
13 : romout=0;
12 : romout=0;
11 : romout=0;
10 : romout=0;
9 : romout=0;
8 : romout=0;
7 : romout=0;
6 : romout=0;
5 : romout=0;
4 : romout=0;
3 : romout=0;
2 : romout=0;
1 : romout=0;
endcase
end
endmodule