module test;
  initial
    begin
      $display("hi");
    end
endmodule

